library verilog;
use verilog.vl_types.all;
entity TB_RAM2 is
end TB_RAM2;
