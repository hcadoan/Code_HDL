library verilog;
use verilog.vl_types.all;
entity TB_baitap7 is
end TB_baitap7;
