library verilog;
use verilog.vl_types.all;
entity TB_RAM1 is
end TB_RAM1;
