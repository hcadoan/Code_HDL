library verilog;
use verilog.vl_types.all;
entity TB_baitap is
end TB_baitap;
