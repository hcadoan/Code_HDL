library verilog;
use verilog.vl_types.all;
entity TB_add4bit is
end TB_add4bit;
