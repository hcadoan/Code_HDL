library verilog;
use verilog.vl_types.all;
entity TB_IC7485 is
end TB_IC7485;
