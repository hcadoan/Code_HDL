library verilog;
use verilog.vl_types.all;
entity TB_RAM_cau2 is
end TB_RAM_cau2;
