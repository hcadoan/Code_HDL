library verilog;
use verilog.vl_types.all;
entity TB_FSM2 is
end TB_FSM2;
