library verilog;
use verilog.vl_types.all;
entity TB_ROM1 is
end TB_ROM1;
