library verilog;
use verilog.vl_types.all;
entity bai4_1 is
    port(
        ck              : in     vl_logic;
        t               : in     vl_logic;
        rs              : in     vl_logic;
        q               : out    vl_logic
    );
end bai4_1;
