library verilog;
use verilog.vl_types.all;
entity TB_nhan4bit is
end TB_nhan4bit;
