library verilog;
use verilog.vl_types.all;
entity TB_mux81_4bit is
end TB_mux81_4bit;
