library verilog;
use verilog.vl_types.all;
entity TB_mux21_8bit is
end TB_mux21_8bit;
