library verilog;
use verilog.vl_types.all;
entity TB_FSM is
end TB_FSM;
