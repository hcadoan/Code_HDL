library verilog;
use verilog.vl_types.all;
entity TB_mux51_led7 is
end TB_mux51_led7;
