library verilog;
use verilog.vl_types.all;
entity fsm1011_vlg_vec_tst is
end fsm1011_vlg_vec_tst;
