library verilog;
use verilog.vl_types.all;
entity TB_demux_18 is
end TB_demux_18;
