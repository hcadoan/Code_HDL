library verilog;
use verilog.vl_types.all;
entity TB_nhan_cong is
end TB_nhan_cong;
