library verilog;
use verilog.vl_types.all;
entity TB_baitap4 is
end TB_baitap4;
