library verilog;
use verilog.vl_types.all;
entity TB_mux51 is
end TB_mux51;
