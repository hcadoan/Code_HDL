library verilog;
use verilog.vl_types.all;
entity TB_nhancong_3bit is
end TB_nhancong_3bit;
