library verilog;
use verilog.vl_types.all;
entity TB_IC74LS151 is
end TB_IC74LS151;
