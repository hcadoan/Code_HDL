library verilog;
use verilog.vl_types.all;
entity mux21_8bit is
    port(
        A               : in     vl_logic_vector(7 downto 0);
        B               : in     vl_logic_vector(7 downto 0);
        S               : in     vl_logic;
        Y               : out    vl_logic_vector(7 downto 0)
    );
end mux21_8bit;
