library verilog;
use verilog.vl_types.all;
entity TB_FSM3 is
end TB_FSM3;
