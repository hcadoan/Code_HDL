library verilog;
use verilog.vl_types.all;
entity TB_bai4_1 is
end TB_bai4_1;
