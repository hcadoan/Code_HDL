library verilog;
use verilog.vl_types.all;
entity bt_vlg_vec_tst is
end bt_vlg_vec_tst;
