library verilog;
use verilog.vl_types.all;
entity cau4_vlg_vec_tst is
end cau4_vlg_vec_tst;
