library verilog;
use verilog.vl_types.all;
entity TB_IC82C19 is
end TB_IC82C19;
