library verilog;
use verilog.vl_types.all;
entity TB_FSM5 is
end TB_FSM5;
