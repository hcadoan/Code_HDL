library verilog;
use verilog.vl_types.all;
entity ss4bit_vlg_vec_tst is
end ss4bit_vlg_vec_tst;
