library verilog;
use verilog.vl_types.all;
entity TB_FSM8 is
end TB_FSM8;
