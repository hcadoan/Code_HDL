library verilog;
use verilog.vl_types.all;
entity TB_bai9 is
end TB_bai9;
