library verilog;
use verilog.vl_types.all;
entity TB_FSM7 is
end TB_FSM7;
