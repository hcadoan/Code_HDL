library verilog;
use verilog.vl_types.all;
entity TB_HAPPY is
end TB_HAPPY;
