library verilog;
use verilog.vl_types.all;
entity TB_demux14_4bit is
end TB_demux14_4bit;
