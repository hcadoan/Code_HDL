library verilog;
use verilog.vl_types.all;
entity TB_bai5_ff is
end TB_bai5_ff;
