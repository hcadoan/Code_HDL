library verilog;
use verilog.vl_types.all;
entity TB_aaa is
end TB_aaa;
