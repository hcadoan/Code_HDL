library verilog;
use verilog.vl_types.all;
entity TB_bt10 is
end TB_bt10;
