library verilog;
use verilog.vl_types.all;
entity TB_FSM9 is
end TB_FSM9;
