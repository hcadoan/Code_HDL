library verilog;
use verilog.vl_types.all;
entity bcd3digit_vlg_vec_tst is
end bcd3digit_vlg_vec_tst;
