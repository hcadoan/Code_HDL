library verilog;
use verilog.vl_types.all;
entity TB_bai2_ram is
end TB_bai2_ram;
