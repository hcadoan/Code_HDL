library verilog;
use verilog.vl_types.all;
entity TB_mux81_8led7 is
end TB_mux81_8led7;
