library verilog;
use verilog.vl_types.all;
entity TB_ROM is
end TB_ROM;
