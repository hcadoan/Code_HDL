library verilog;
use verilog.vl_types.all;
entity TB_RAM is
end TB_RAM;
