library verilog;
use verilog.vl_types.all;
entity TB_baitap2 is
end TB_baitap2;
