library verilog;
use verilog.vl_types.all;
entity cau3_vlg_vec_tst is
end cau3_vlg_vec_tst;
