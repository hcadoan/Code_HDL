library verilog;
use verilog.vl_types.all;
entity TB_add8bit is
end TB_add8bit;
