library verilog;
use verilog.vl_types.all;
entity TB_FSM_cau3 is
end TB_FSM_cau3;
