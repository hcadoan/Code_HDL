library verilog;
use verilog.vl_types.all;
entity TB_baitap3 is
end TB_baitap3;
