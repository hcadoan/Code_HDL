library verilog;
use verilog.vl_types.all;
entity nhan4bit_vlg_vec_tst is
end nhan4bit_vlg_vec_tst;
