library verilog;
use verilog.vl_types.all;
entity TB_ROM_cau1 is
end TB_ROM_cau1;
