library verilog;
use verilog.vl_types.all;
entity bcd_mod60_vlg_vec_tst is
end bcd_mod60_vlg_vec_tst;
